library verilog;
use verilog.vl_types.all;
entity ten_counter_vlg_vec_tst is
end ten_counter_vlg_vec_tst;
