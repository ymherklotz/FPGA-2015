library verilog;
use verilog.vl_types.all;
entity bcd_to_display_vlg_vec_tst is
end bcd_to_display_vlg_vec_tst;
